module and_module(a, b, o);
  input a;
  input b;
  output o;
  wire a, b, o;
  assign o = a & b;
endmodule
